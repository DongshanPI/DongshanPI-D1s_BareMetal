
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h4f542320;
    ram_cell[       1] = 32'h0;  // 32'he576fe62;
    ram_cell[       2] = 32'h0;  // 32'h75241a41;
    ram_cell[       3] = 32'h0;  // 32'h4f48d574;
    ram_cell[       4] = 32'h0;  // 32'h7a4687f3;
    ram_cell[       5] = 32'h0;  // 32'h9e298cb0;
    ram_cell[       6] = 32'h0;  // 32'hbad5c319;
    ram_cell[       7] = 32'h0;  // 32'h5c340c71;
    ram_cell[       8] = 32'h0;  // 32'h116d5889;
    ram_cell[       9] = 32'h0;  // 32'ha9eea31e;
    ram_cell[      10] = 32'h0;  // 32'h94f53a16;
    ram_cell[      11] = 32'h0;  // 32'hcee93bc9;
    ram_cell[      12] = 32'h0;  // 32'hb9f52b12;
    ram_cell[      13] = 32'h0;  // 32'hc618d382;
    ram_cell[      14] = 32'h0;  // 32'h4c515451;
    ram_cell[      15] = 32'h0;  // 32'h79c58b5e;
    ram_cell[      16] = 32'h0;  // 32'h4ec66b3f;
    ram_cell[      17] = 32'h0;  // 32'h5c420c25;
    ram_cell[      18] = 32'h0;  // 32'h140676f0;
    ram_cell[      19] = 32'h0;  // 32'h77c0fd42;
    ram_cell[      20] = 32'h0;  // 32'ha866e26f;
    ram_cell[      21] = 32'h0;  // 32'hc6fb7d00;
    ram_cell[      22] = 32'h0;  // 32'h92db61ad;
    ram_cell[      23] = 32'h0;  // 32'hf8fbaab4;
    ram_cell[      24] = 32'h0;  // 32'h2bb94160;
    ram_cell[      25] = 32'h0;  // 32'h2db8062a;
    ram_cell[      26] = 32'h0;  // 32'hc6cd4ef2;
    ram_cell[      27] = 32'h0;  // 32'hd9a0fcf4;
    ram_cell[      28] = 32'h0;  // 32'h36d1de19;
    ram_cell[      29] = 32'h0;  // 32'h637f4ce8;
    ram_cell[      30] = 32'h0;  // 32'h5d1ba96f;
    ram_cell[      31] = 32'h0;  // 32'hfb908b1e;
    ram_cell[      32] = 32'h0;  // 32'h25db44b3;
    ram_cell[      33] = 32'h0;  // 32'hbecfcbbf;
    ram_cell[      34] = 32'h0;  // 32'h5df516e2;
    ram_cell[      35] = 32'h0;  // 32'hc926042e;
    ram_cell[      36] = 32'h0;  // 32'h03f2140f;
    ram_cell[      37] = 32'h0;  // 32'ha897b4eb;
    ram_cell[      38] = 32'h0;  // 32'h50922263;
    ram_cell[      39] = 32'h0;  // 32'h02b914dc;
    ram_cell[      40] = 32'h0;  // 32'hef54290b;
    ram_cell[      41] = 32'h0;  // 32'h19920a80;
    ram_cell[      42] = 32'h0;  // 32'hc3fdb6fa;
    ram_cell[      43] = 32'h0;  // 32'hffc45d84;
    ram_cell[      44] = 32'h0;  // 32'h81285860;
    ram_cell[      45] = 32'h0;  // 32'h4e057836;
    ram_cell[      46] = 32'h0;  // 32'hf5ab864a;
    ram_cell[      47] = 32'h0;  // 32'h6cde453f;
    ram_cell[      48] = 32'h0;  // 32'h3c39905e;
    ram_cell[      49] = 32'h0;  // 32'h84e3e2ce;
    ram_cell[      50] = 32'h0;  // 32'h06b18028;
    ram_cell[      51] = 32'h0;  // 32'he79aa241;
    ram_cell[      52] = 32'h0;  // 32'h08fb80de;
    ram_cell[      53] = 32'h0;  // 32'he7b0ede9;
    ram_cell[      54] = 32'h0;  // 32'h3e697ca3;
    ram_cell[      55] = 32'h0;  // 32'ha3e93015;
    ram_cell[      56] = 32'h0;  // 32'h3e3f64df;
    ram_cell[      57] = 32'h0;  // 32'h3f110810;
    ram_cell[      58] = 32'h0;  // 32'h27d43890;
    ram_cell[      59] = 32'h0;  // 32'h004e40ae;
    ram_cell[      60] = 32'h0;  // 32'hb4ebbb86;
    ram_cell[      61] = 32'h0;  // 32'ha5d466e7;
    ram_cell[      62] = 32'h0;  // 32'hd53b55b8;
    ram_cell[      63] = 32'h0;  // 32'hfc67661a;
    ram_cell[      64] = 32'h0;  // 32'ha73b0e2a;
    ram_cell[      65] = 32'h0;  // 32'ha732260b;
    ram_cell[      66] = 32'h0;  // 32'h2bd4950e;
    ram_cell[      67] = 32'h0;  // 32'haa30a5e9;
    ram_cell[      68] = 32'h0;  // 32'hb37cb060;
    ram_cell[      69] = 32'h0;  // 32'haedf35a5;
    ram_cell[      70] = 32'h0;  // 32'h4bb887c1;
    ram_cell[      71] = 32'h0;  // 32'h7fa18578;
    ram_cell[      72] = 32'h0;  // 32'h19bcc264;
    ram_cell[      73] = 32'h0;  // 32'h3a6c3a41;
    ram_cell[      74] = 32'h0;  // 32'h70b4b9ab;
    ram_cell[      75] = 32'h0;  // 32'h2f96e138;
    ram_cell[      76] = 32'h0;  // 32'h0cc566ce;
    ram_cell[      77] = 32'h0;  // 32'he11d39c5;
    ram_cell[      78] = 32'h0;  // 32'ha3b48ffe;
    ram_cell[      79] = 32'h0;  // 32'h86c38af8;
    ram_cell[      80] = 32'h0;  // 32'h971308df;
    ram_cell[      81] = 32'h0;  // 32'he624a236;
    ram_cell[      82] = 32'h0;  // 32'h6d1c2d8d;
    ram_cell[      83] = 32'h0;  // 32'h8b89435a;
    ram_cell[      84] = 32'h0;  // 32'h383458f7;
    ram_cell[      85] = 32'h0;  // 32'h8d2555b2;
    ram_cell[      86] = 32'h0;  // 32'hba5a3362;
    ram_cell[      87] = 32'h0;  // 32'h495e5636;
    ram_cell[      88] = 32'h0;  // 32'h3cd60982;
    ram_cell[      89] = 32'h0;  // 32'h2dadd57b;
    ram_cell[      90] = 32'h0;  // 32'h926836f1;
    ram_cell[      91] = 32'h0;  // 32'h26eeb980;
    ram_cell[      92] = 32'h0;  // 32'h4d72b4b4;
    ram_cell[      93] = 32'h0;  // 32'hfe3eae42;
    ram_cell[      94] = 32'h0;  // 32'he96a685c;
    ram_cell[      95] = 32'h0;  // 32'ha5749fa4;
    ram_cell[      96] = 32'h0;  // 32'h8b812c00;
    ram_cell[      97] = 32'h0;  // 32'h1e495ac7;
    ram_cell[      98] = 32'h0;  // 32'hc5e19d30;
    ram_cell[      99] = 32'h0;  // 32'h5ff32665;
    ram_cell[     100] = 32'h0;  // 32'h9f9215f1;
    ram_cell[     101] = 32'h0;  // 32'he02cfa0d;
    ram_cell[     102] = 32'h0;  // 32'ha2894b96;
    ram_cell[     103] = 32'h0;  // 32'h047492e6;
    ram_cell[     104] = 32'h0;  // 32'hf0734038;
    ram_cell[     105] = 32'h0;  // 32'hd8b2fae9;
    ram_cell[     106] = 32'h0;  // 32'h68fa47da;
    ram_cell[     107] = 32'h0;  // 32'h03223602;
    ram_cell[     108] = 32'h0;  // 32'h25c21ede;
    ram_cell[     109] = 32'h0;  // 32'h82c8a81f;
    ram_cell[     110] = 32'h0;  // 32'h1b1eee0e;
    ram_cell[     111] = 32'h0;  // 32'hd29be268;
    ram_cell[     112] = 32'h0;  // 32'hca237fdb;
    ram_cell[     113] = 32'h0;  // 32'h2f35dbce;
    ram_cell[     114] = 32'h0;  // 32'hb23017fe;
    ram_cell[     115] = 32'h0;  // 32'h5f97a387;
    ram_cell[     116] = 32'h0;  // 32'h65ce4d51;
    ram_cell[     117] = 32'h0;  // 32'h7160f348;
    ram_cell[     118] = 32'h0;  // 32'h6b2a2605;
    ram_cell[     119] = 32'h0;  // 32'h38341369;
    ram_cell[     120] = 32'h0;  // 32'he1679efa;
    ram_cell[     121] = 32'h0;  // 32'h22234e74;
    ram_cell[     122] = 32'h0;  // 32'h406740c7;
    ram_cell[     123] = 32'h0;  // 32'hea6f226b;
    ram_cell[     124] = 32'h0;  // 32'hefa0bbb1;
    ram_cell[     125] = 32'h0;  // 32'h925ba4fd;
    ram_cell[     126] = 32'h0;  // 32'h77d09537;
    ram_cell[     127] = 32'h0;  // 32'h2ea77a61;
    ram_cell[     128] = 32'h0;  // 32'h353fd766;
    ram_cell[     129] = 32'h0;  // 32'hfa96cc15;
    ram_cell[     130] = 32'h0;  // 32'hcec7a6b3;
    ram_cell[     131] = 32'h0;  // 32'h10d58775;
    ram_cell[     132] = 32'h0;  // 32'hd8e6a962;
    ram_cell[     133] = 32'h0;  // 32'h03e4c9f5;
    ram_cell[     134] = 32'h0;  // 32'h40e787fa;
    ram_cell[     135] = 32'h0;  // 32'h070e5ee6;
    ram_cell[     136] = 32'h0;  // 32'h5bac6e49;
    ram_cell[     137] = 32'h0;  // 32'h07b2528c;
    ram_cell[     138] = 32'h0;  // 32'h4109d9cc;
    ram_cell[     139] = 32'h0;  // 32'he7cad4df;
    ram_cell[     140] = 32'h0;  // 32'hb138a485;
    ram_cell[     141] = 32'h0;  // 32'h86d51760;
    ram_cell[     142] = 32'h0;  // 32'hf0ef0df5;
    ram_cell[     143] = 32'h0;  // 32'h007b2c74;
    ram_cell[     144] = 32'h0;  // 32'h9e3277a2;
    ram_cell[     145] = 32'h0;  // 32'h1abcbd90;
    ram_cell[     146] = 32'h0;  // 32'h93d1f79f;
    ram_cell[     147] = 32'h0;  // 32'hc29534b1;
    ram_cell[     148] = 32'h0;  // 32'ha994cebb;
    ram_cell[     149] = 32'h0;  // 32'h2ede5a36;
    ram_cell[     150] = 32'h0;  // 32'hdac67121;
    ram_cell[     151] = 32'h0;  // 32'hf3c65633;
    ram_cell[     152] = 32'h0;  // 32'hbf2842e6;
    ram_cell[     153] = 32'h0;  // 32'hb64a510e;
    ram_cell[     154] = 32'h0;  // 32'h0d191a56;
    ram_cell[     155] = 32'h0;  // 32'h39e933df;
    ram_cell[     156] = 32'h0;  // 32'h56379c7b;
    ram_cell[     157] = 32'h0;  // 32'hf870dbc1;
    ram_cell[     158] = 32'h0;  // 32'hd7cdb899;
    ram_cell[     159] = 32'h0;  // 32'h45e24a2e;
    ram_cell[     160] = 32'h0;  // 32'ha4bf5628;
    ram_cell[     161] = 32'h0;  // 32'h6d0e5f61;
    ram_cell[     162] = 32'h0;  // 32'h9318d51c;
    ram_cell[     163] = 32'h0;  // 32'h90b5ab19;
    ram_cell[     164] = 32'h0;  // 32'h65a4be01;
    ram_cell[     165] = 32'h0;  // 32'h9fab1b4c;
    ram_cell[     166] = 32'h0;  // 32'he087721d;
    ram_cell[     167] = 32'h0;  // 32'hb6c68ad2;
    ram_cell[     168] = 32'h0;  // 32'h7944e68e;
    ram_cell[     169] = 32'h0;  // 32'hc7878fc2;
    ram_cell[     170] = 32'h0;  // 32'h0c8ca70e;
    ram_cell[     171] = 32'h0;  // 32'h4e005b72;
    ram_cell[     172] = 32'h0;  // 32'hc3f8ba60;
    ram_cell[     173] = 32'h0;  // 32'h4c3814d2;
    ram_cell[     174] = 32'h0;  // 32'h276e9c4b;
    ram_cell[     175] = 32'h0;  // 32'h3df4b1da;
    ram_cell[     176] = 32'h0;  // 32'h69a6d3bc;
    ram_cell[     177] = 32'h0;  // 32'hc148ae43;
    ram_cell[     178] = 32'h0;  // 32'h5994312e;
    ram_cell[     179] = 32'h0;  // 32'ha21d88b1;
    ram_cell[     180] = 32'h0;  // 32'ha24f2857;
    ram_cell[     181] = 32'h0;  // 32'h6602a295;
    ram_cell[     182] = 32'h0;  // 32'h487f1d93;
    ram_cell[     183] = 32'h0;  // 32'h76ab194c;
    ram_cell[     184] = 32'h0;  // 32'hacc214db;
    ram_cell[     185] = 32'h0;  // 32'hbd90a3f6;
    ram_cell[     186] = 32'h0;  // 32'h479ad9db;
    ram_cell[     187] = 32'h0;  // 32'h676f5418;
    ram_cell[     188] = 32'h0;  // 32'h81551936;
    ram_cell[     189] = 32'h0;  // 32'h23619575;
    ram_cell[     190] = 32'h0;  // 32'hb0e231b2;
    ram_cell[     191] = 32'h0;  // 32'h7e7a787c;
    ram_cell[     192] = 32'h0;  // 32'h075354df;
    ram_cell[     193] = 32'h0;  // 32'h99e1f6dd;
    ram_cell[     194] = 32'h0;  // 32'h07156877;
    ram_cell[     195] = 32'h0;  // 32'h4716a05d;
    ram_cell[     196] = 32'h0;  // 32'h58513ed1;
    ram_cell[     197] = 32'h0;  // 32'h78b3b4ca;
    ram_cell[     198] = 32'h0;  // 32'h70300ad8;
    ram_cell[     199] = 32'h0;  // 32'h19c2aae7;
    ram_cell[     200] = 32'h0;  // 32'h179ae2c0;
    ram_cell[     201] = 32'h0;  // 32'h527b6083;
    ram_cell[     202] = 32'h0;  // 32'h779ed944;
    ram_cell[     203] = 32'h0;  // 32'h3915b626;
    ram_cell[     204] = 32'h0;  // 32'hf98049ab;
    ram_cell[     205] = 32'h0;  // 32'h5d7549c7;
    ram_cell[     206] = 32'h0;  // 32'h1f337b9f;
    ram_cell[     207] = 32'h0;  // 32'hbc6e2d89;
    ram_cell[     208] = 32'h0;  // 32'hda98b4f9;
    ram_cell[     209] = 32'h0;  // 32'h0ca14530;
    ram_cell[     210] = 32'h0;  // 32'h19d3521a;
    ram_cell[     211] = 32'h0;  // 32'hdd7fc744;
    ram_cell[     212] = 32'h0;  // 32'hd9497930;
    ram_cell[     213] = 32'h0;  // 32'ha951f730;
    ram_cell[     214] = 32'h0;  // 32'h1a485d44;
    ram_cell[     215] = 32'h0;  // 32'h5892b3c2;
    ram_cell[     216] = 32'h0;  // 32'hc2d42a94;
    ram_cell[     217] = 32'h0;  // 32'hd2ac199f;
    ram_cell[     218] = 32'h0;  // 32'hefef79d5;
    ram_cell[     219] = 32'h0;  // 32'hdf0cc79c;
    ram_cell[     220] = 32'h0;  // 32'hade655a1;
    ram_cell[     221] = 32'h0;  // 32'h32c7899b;
    ram_cell[     222] = 32'h0;  // 32'h183f276f;
    ram_cell[     223] = 32'h0;  // 32'h8554ce8d;
    ram_cell[     224] = 32'h0;  // 32'h2aef18e2;
    ram_cell[     225] = 32'h0;  // 32'h5a0e6953;
    ram_cell[     226] = 32'h0;  // 32'h4c243020;
    ram_cell[     227] = 32'h0;  // 32'h7ba463e6;
    ram_cell[     228] = 32'h0;  // 32'hbe68fcb9;
    ram_cell[     229] = 32'h0;  // 32'ha93eb87b;
    ram_cell[     230] = 32'h0;  // 32'h7a3ceeff;
    ram_cell[     231] = 32'h0;  // 32'h912493e9;
    ram_cell[     232] = 32'h0;  // 32'h35e64cfb;
    ram_cell[     233] = 32'h0;  // 32'ha8e86e7c;
    ram_cell[     234] = 32'h0;  // 32'h0d0997de;
    ram_cell[     235] = 32'h0;  // 32'h9f7a5631;
    ram_cell[     236] = 32'h0;  // 32'h8f0148ec;
    ram_cell[     237] = 32'h0;  // 32'hfebf1cd3;
    ram_cell[     238] = 32'h0;  // 32'h3f856cd4;
    ram_cell[     239] = 32'h0;  // 32'h6091f711;
    ram_cell[     240] = 32'h0;  // 32'h3584bd41;
    ram_cell[     241] = 32'h0;  // 32'h3600190d;
    ram_cell[     242] = 32'h0;  // 32'h82d66b85;
    ram_cell[     243] = 32'h0;  // 32'h7b75b906;
    ram_cell[     244] = 32'h0;  // 32'h0a6fc712;
    ram_cell[     245] = 32'h0;  // 32'h7e693836;
    ram_cell[     246] = 32'h0;  // 32'hfd4a0441;
    ram_cell[     247] = 32'h0;  // 32'h7fbd4d37;
    ram_cell[     248] = 32'h0;  // 32'h258db53c;
    ram_cell[     249] = 32'h0;  // 32'h514d77b5;
    ram_cell[     250] = 32'h0;  // 32'hc95fdc42;
    ram_cell[     251] = 32'h0;  // 32'hba8e15ba;
    ram_cell[     252] = 32'h0;  // 32'hffe6f889;
    ram_cell[     253] = 32'h0;  // 32'h6329e0c9;
    ram_cell[     254] = 32'h0;  // 32'h60749cab;
    ram_cell[     255] = 32'h0;  // 32'hf5d41d5b;
    // src matrix A
    ram_cell[     256] = 32'h34802979;
    ram_cell[     257] = 32'hf5ea385f;
    ram_cell[     258] = 32'hc21e78a7;
    ram_cell[     259] = 32'h4f8d63d4;
    ram_cell[     260] = 32'h5059d3f5;
    ram_cell[     261] = 32'he95c07e9;
    ram_cell[     262] = 32'hc0767230;
    ram_cell[     263] = 32'h127078a4;
    ram_cell[     264] = 32'h8c251245;
    ram_cell[     265] = 32'h84d24fdd;
    ram_cell[     266] = 32'ha63629f0;
    ram_cell[     267] = 32'h344846e7;
    ram_cell[     268] = 32'hf40f11e2;
    ram_cell[     269] = 32'h9eb21e36;
    ram_cell[     270] = 32'h93e4fbb3;
    ram_cell[     271] = 32'h9b8d2efb;
    ram_cell[     272] = 32'hae50fa1d;
    ram_cell[     273] = 32'hecadc2db;
    ram_cell[     274] = 32'h3cab352a;
    ram_cell[     275] = 32'hca85010e;
    ram_cell[     276] = 32'h9b88f719;
    ram_cell[     277] = 32'h58c17235;
    ram_cell[     278] = 32'h2f8a98ca;
    ram_cell[     279] = 32'h1362d566;
    ram_cell[     280] = 32'hc2347f5a;
    ram_cell[     281] = 32'h18b3c0fe;
    ram_cell[     282] = 32'h1c9b0f4c;
    ram_cell[     283] = 32'h7b709d43;
    ram_cell[     284] = 32'h8a4f9eb6;
    ram_cell[     285] = 32'h8e4c8540;
    ram_cell[     286] = 32'he399d889;
    ram_cell[     287] = 32'hca364286;
    ram_cell[     288] = 32'hee94c150;
    ram_cell[     289] = 32'h9513b0a0;
    ram_cell[     290] = 32'h9f9d13c3;
    ram_cell[     291] = 32'h098fd433;
    ram_cell[     292] = 32'hc6d74e37;
    ram_cell[     293] = 32'h1dc00c81;
    ram_cell[     294] = 32'hc6d755c9;
    ram_cell[     295] = 32'ha4b6678c;
    ram_cell[     296] = 32'he0739216;
    ram_cell[     297] = 32'h4b740934;
    ram_cell[     298] = 32'h2cde455a;
    ram_cell[     299] = 32'h055617ae;
    ram_cell[     300] = 32'hb859eedf;
    ram_cell[     301] = 32'hdc8f85ca;
    ram_cell[     302] = 32'h6b68e832;
    ram_cell[     303] = 32'h098d4d2a;
    ram_cell[     304] = 32'h7784e913;
    ram_cell[     305] = 32'h12db286b;
    ram_cell[     306] = 32'h00acce46;
    ram_cell[     307] = 32'h00e8fbb7;
    ram_cell[     308] = 32'hbfbbfed2;
    ram_cell[     309] = 32'h9dea31f2;
    ram_cell[     310] = 32'h3eb1dc40;
    ram_cell[     311] = 32'h49dfefc0;
    ram_cell[     312] = 32'hfecd0811;
    ram_cell[     313] = 32'hf28e8110;
    ram_cell[     314] = 32'hfc57750e;
    ram_cell[     315] = 32'hd034fca4;
    ram_cell[     316] = 32'h2feebed4;
    ram_cell[     317] = 32'h1c652425;
    ram_cell[     318] = 32'he0997154;
    ram_cell[     319] = 32'h2a70c8c8;
    ram_cell[     320] = 32'h3a34b748;
    ram_cell[     321] = 32'ha0b343e4;
    ram_cell[     322] = 32'ha2caebc8;
    ram_cell[     323] = 32'h8e529268;
    ram_cell[     324] = 32'h7decb6b1;
    ram_cell[     325] = 32'h10003965;
    ram_cell[     326] = 32'h1945f3a0;
    ram_cell[     327] = 32'hc38ece9f;
    ram_cell[     328] = 32'h15d6eeba;
    ram_cell[     329] = 32'h18beca0d;
    ram_cell[     330] = 32'h1d6852ca;
    ram_cell[     331] = 32'h1f0e4d2c;
    ram_cell[     332] = 32'ha15ec55c;
    ram_cell[     333] = 32'hd3a89350;
    ram_cell[     334] = 32'h1c5c8cba;
    ram_cell[     335] = 32'hca36d3f1;
    ram_cell[     336] = 32'haa354111;
    ram_cell[     337] = 32'h2bde03ab;
    ram_cell[     338] = 32'h310d1e3a;
    ram_cell[     339] = 32'h3501a6ca;
    ram_cell[     340] = 32'h450851f5;
    ram_cell[     341] = 32'h64d4982b;
    ram_cell[     342] = 32'h4b2e26d1;
    ram_cell[     343] = 32'hcd0be3c6;
    ram_cell[     344] = 32'h48eea40b;
    ram_cell[     345] = 32'h29527e09;
    ram_cell[     346] = 32'hd44ffa94;
    ram_cell[     347] = 32'hce86fb39;
    ram_cell[     348] = 32'hec8d688b;
    ram_cell[     349] = 32'h3596c407;
    ram_cell[     350] = 32'h3bc668e1;
    ram_cell[     351] = 32'hfc341f32;
    ram_cell[     352] = 32'hd21efd98;
    ram_cell[     353] = 32'h7266f3af;
    ram_cell[     354] = 32'hde4e3805;
    ram_cell[     355] = 32'hf856a03f;
    ram_cell[     356] = 32'h52c222c7;
    ram_cell[     357] = 32'h4c12b9ba;
    ram_cell[     358] = 32'h9efa4237;
    ram_cell[     359] = 32'h5fbcbf09;
    ram_cell[     360] = 32'hb9fce6b2;
    ram_cell[     361] = 32'h37d95eaf;
    ram_cell[     362] = 32'hd6fb9d67;
    ram_cell[     363] = 32'ha1bbfbf0;
    ram_cell[     364] = 32'h35bd79f3;
    ram_cell[     365] = 32'h38f7deae;
    ram_cell[     366] = 32'hf1f8e1fa;
    ram_cell[     367] = 32'h9e84654b;
    ram_cell[     368] = 32'h0d487e49;
    ram_cell[     369] = 32'hbecc6697;
    ram_cell[     370] = 32'hb19c8266;
    ram_cell[     371] = 32'h2d6e6fe5;
    ram_cell[     372] = 32'h3a224912;
    ram_cell[     373] = 32'h56a5bbe5;
    ram_cell[     374] = 32'hc5c8d159;
    ram_cell[     375] = 32'h990b1682;
    ram_cell[     376] = 32'h779ee895;
    ram_cell[     377] = 32'hc8b21e8f;
    ram_cell[     378] = 32'h8d0dfe29;
    ram_cell[     379] = 32'hb4fec42f;
    ram_cell[     380] = 32'hf043eb29;
    ram_cell[     381] = 32'hdc12b7ce;
    ram_cell[     382] = 32'haa198c53;
    ram_cell[     383] = 32'h51cf9a85;
    ram_cell[     384] = 32'hb2778727;
    ram_cell[     385] = 32'hee5870bc;
    ram_cell[     386] = 32'h48b29b2e;
    ram_cell[     387] = 32'hbf843f52;
    ram_cell[     388] = 32'h9ff10d96;
    ram_cell[     389] = 32'h4b79ea84;
    ram_cell[     390] = 32'hf1ca2f5a;
    ram_cell[     391] = 32'hf5e96481;
    ram_cell[     392] = 32'h9ced6638;
    ram_cell[     393] = 32'h9c2514be;
    ram_cell[     394] = 32'h474464b7;
    ram_cell[     395] = 32'hfaf1db5c;
    ram_cell[     396] = 32'hda8f2c8f;
    ram_cell[     397] = 32'h9a8506fa;
    ram_cell[     398] = 32'h796b8492;
    ram_cell[     399] = 32'h73fcdc61;
    ram_cell[     400] = 32'h7f868a38;
    ram_cell[     401] = 32'h8d375dc0;
    ram_cell[     402] = 32'hd29c9d07;
    ram_cell[     403] = 32'h7cb3ac3f;
    ram_cell[     404] = 32'h47b23478;
    ram_cell[     405] = 32'h89aa3c5f;
    ram_cell[     406] = 32'hc2d8dbc4;
    ram_cell[     407] = 32'h6210f969;
    ram_cell[     408] = 32'h05540701;
    ram_cell[     409] = 32'ha70f4574;
    ram_cell[     410] = 32'h57a8dea1;
    ram_cell[     411] = 32'h76a487f2;
    ram_cell[     412] = 32'hdb789d95;
    ram_cell[     413] = 32'h4fc9cb14;
    ram_cell[     414] = 32'hebc87c4b;
    ram_cell[     415] = 32'ha74fcda8;
    ram_cell[     416] = 32'h03111971;
    ram_cell[     417] = 32'h2ccb46c3;
    ram_cell[     418] = 32'h6819f77a;
    ram_cell[     419] = 32'hbd198f5b;
    ram_cell[     420] = 32'h6678dcde;
    ram_cell[     421] = 32'h3917762a;
    ram_cell[     422] = 32'h0d6bdae3;
    ram_cell[     423] = 32'h7433d774;
    ram_cell[     424] = 32'hec7bd607;
    ram_cell[     425] = 32'hde96749e;
    ram_cell[     426] = 32'hd18ce89a;
    ram_cell[     427] = 32'h916d1415;
    ram_cell[     428] = 32'h4fabde3a;
    ram_cell[     429] = 32'he68cb6a5;
    ram_cell[     430] = 32'h236ee634;
    ram_cell[     431] = 32'hcec3e277;
    ram_cell[     432] = 32'hee60ce28;
    ram_cell[     433] = 32'h7ede246e;
    ram_cell[     434] = 32'h3cfadd32;
    ram_cell[     435] = 32'h919febc4;
    ram_cell[     436] = 32'hecad1191;
    ram_cell[     437] = 32'h9caa1505;
    ram_cell[     438] = 32'h6fc83f5c;
    ram_cell[     439] = 32'hd46f7844;
    ram_cell[     440] = 32'h5294eb32;
    ram_cell[     441] = 32'h221389ea;
    ram_cell[     442] = 32'h4a4d8983;
    ram_cell[     443] = 32'he0f8067d;
    ram_cell[     444] = 32'h3c5b6e9d;
    ram_cell[     445] = 32'h17d8709d;
    ram_cell[     446] = 32'hc6a94775;
    ram_cell[     447] = 32'h9995486f;
    ram_cell[     448] = 32'hff184be8;
    ram_cell[     449] = 32'h25f9b2cb;
    ram_cell[     450] = 32'h465a5ba3;
    ram_cell[     451] = 32'h8458852b;
    ram_cell[     452] = 32'hdcfc7645;
    ram_cell[     453] = 32'hf996f22c;
    ram_cell[     454] = 32'h8f6c360f;
    ram_cell[     455] = 32'h65aee623;
    ram_cell[     456] = 32'hc9d958e7;
    ram_cell[     457] = 32'h00ffa61d;
    ram_cell[     458] = 32'hc2f85d15;
    ram_cell[     459] = 32'hd511baf2;
    ram_cell[     460] = 32'h6755968a;
    ram_cell[     461] = 32'h1fbc29c0;
    ram_cell[     462] = 32'hf3072831;
    ram_cell[     463] = 32'h5f5f0bbc;
    ram_cell[     464] = 32'he92be7d5;
    ram_cell[     465] = 32'hafa8e34f;
    ram_cell[     466] = 32'hdd9f20e9;
    ram_cell[     467] = 32'hddecddd9;
    ram_cell[     468] = 32'h42df489b;
    ram_cell[     469] = 32'hc0348d43;
    ram_cell[     470] = 32'h6b0372cd;
    ram_cell[     471] = 32'hfbf50607;
    ram_cell[     472] = 32'h30f6d853;
    ram_cell[     473] = 32'hd2736431;
    ram_cell[     474] = 32'haaf57b19;
    ram_cell[     475] = 32'h2d2810e5;
    ram_cell[     476] = 32'h6eacc05f;
    ram_cell[     477] = 32'h50480710;
    ram_cell[     478] = 32'h0250203e;
    ram_cell[     479] = 32'h9c0c4eed;
    ram_cell[     480] = 32'he0e14e38;
    ram_cell[     481] = 32'h2fe441c9;
    ram_cell[     482] = 32'ha0d6aeca;
    ram_cell[     483] = 32'h4b5d0f6d;
    ram_cell[     484] = 32'h2957fb13;
    ram_cell[     485] = 32'haa35dccb;
    ram_cell[     486] = 32'h54b578c9;
    ram_cell[     487] = 32'haf7653b3;
    ram_cell[     488] = 32'h77e83066;
    ram_cell[     489] = 32'h24c5f378;
    ram_cell[     490] = 32'h4c55c5e4;
    ram_cell[     491] = 32'h7e3b69b5;
    ram_cell[     492] = 32'he79d06ba;
    ram_cell[     493] = 32'h471633e3;
    ram_cell[     494] = 32'h1378e714;
    ram_cell[     495] = 32'h1c641d9d;
    ram_cell[     496] = 32'h5f01fd6d;
    ram_cell[     497] = 32'h39f7cc8b;
    ram_cell[     498] = 32'h0f9677d6;
    ram_cell[     499] = 32'h2f504489;
    ram_cell[     500] = 32'h1c5c0ce6;
    ram_cell[     501] = 32'ha1fbdfcf;
    ram_cell[     502] = 32'h8a2946de;
    ram_cell[     503] = 32'h59cabac4;
    ram_cell[     504] = 32'h197d101f;
    ram_cell[     505] = 32'h31c94861;
    ram_cell[     506] = 32'h4796fe47;
    ram_cell[     507] = 32'h1eb2a43d;
    ram_cell[     508] = 32'ha5d6349a;
    ram_cell[     509] = 32'hd2e5f7ce;
    ram_cell[     510] = 32'h3414659d;
    ram_cell[     511] = 32'h3933c9d8;
    // src matrix B
    ram_cell[     512] = 32'hfdd2ccf6;
    ram_cell[     513] = 32'he535905d;
    ram_cell[     514] = 32'ha733ceb0;
    ram_cell[     515] = 32'ha00fc0bd;
    ram_cell[     516] = 32'h9404dc68;
    ram_cell[     517] = 32'h7a8bf7f7;
    ram_cell[     518] = 32'hdfb7a7f0;
    ram_cell[     519] = 32'hed493033;
    ram_cell[     520] = 32'h37a62a17;
    ram_cell[     521] = 32'had8ef068;
    ram_cell[     522] = 32'h7bfeb45a;
    ram_cell[     523] = 32'hcc62c287;
    ram_cell[     524] = 32'h9e4026f1;
    ram_cell[     525] = 32'hd0e7b94c;
    ram_cell[     526] = 32'h31d65aca;
    ram_cell[     527] = 32'h354b70b8;
    ram_cell[     528] = 32'h33584afb;
    ram_cell[     529] = 32'he736ff46;
    ram_cell[     530] = 32'ha30ac32b;
    ram_cell[     531] = 32'h99932bed;
    ram_cell[     532] = 32'h60fafb1f;
    ram_cell[     533] = 32'h88572860;
    ram_cell[     534] = 32'hdbd06f3b;
    ram_cell[     535] = 32'h44a61cfc;
    ram_cell[     536] = 32'h19394a6d;
    ram_cell[     537] = 32'h5efe455b;
    ram_cell[     538] = 32'hcd536a5c;
    ram_cell[     539] = 32'h861d791c;
    ram_cell[     540] = 32'h48e1306b;
    ram_cell[     541] = 32'hdb48add1;
    ram_cell[     542] = 32'hfb4ea412;
    ram_cell[     543] = 32'he141ff94;
    ram_cell[     544] = 32'h5c67aae9;
    ram_cell[     545] = 32'h7d153967;
    ram_cell[     546] = 32'ha365584b;
    ram_cell[     547] = 32'h2fd3d12f;
    ram_cell[     548] = 32'h8fc1844e;
    ram_cell[     549] = 32'h2b6d575b;
    ram_cell[     550] = 32'hd593399f;
    ram_cell[     551] = 32'hc5b5d06d;
    ram_cell[     552] = 32'h7d79d953;
    ram_cell[     553] = 32'h4c2e49a5;
    ram_cell[     554] = 32'ha6ef77af;
    ram_cell[     555] = 32'h8ed10a15;
    ram_cell[     556] = 32'ha4c90260;
    ram_cell[     557] = 32'h19b463f2;
    ram_cell[     558] = 32'h2402486d;
    ram_cell[     559] = 32'h616f115b;
    ram_cell[     560] = 32'h13f47649;
    ram_cell[     561] = 32'hf9989727;
    ram_cell[     562] = 32'hcb79bb3b;
    ram_cell[     563] = 32'hbf30d4a8;
    ram_cell[     564] = 32'h8319bcf0;
    ram_cell[     565] = 32'ha317efc8;
    ram_cell[     566] = 32'h23035491;
    ram_cell[     567] = 32'h34fb48a4;
    ram_cell[     568] = 32'hc87ae36c;
    ram_cell[     569] = 32'he396ccbd;
    ram_cell[     570] = 32'h4516356d;
    ram_cell[     571] = 32'hf3a59620;
    ram_cell[     572] = 32'h89cbc120;
    ram_cell[     573] = 32'h2f10da99;
    ram_cell[     574] = 32'h1c863d6f;
    ram_cell[     575] = 32'h204f5f16;
    ram_cell[     576] = 32'hd5d05868;
    ram_cell[     577] = 32'h5827a6fa;
    ram_cell[     578] = 32'hadb94b66;
    ram_cell[     579] = 32'hf9a5f38b;
    ram_cell[     580] = 32'h9ef4eac4;
    ram_cell[     581] = 32'hf20d871e;
    ram_cell[     582] = 32'h552f9aac;
    ram_cell[     583] = 32'h34fbe673;
    ram_cell[     584] = 32'hba52982c;
    ram_cell[     585] = 32'h868efc4e;
    ram_cell[     586] = 32'hdd29b35b;
    ram_cell[     587] = 32'h68724b24;
    ram_cell[     588] = 32'h4a544bed;
    ram_cell[     589] = 32'h831c435a;
    ram_cell[     590] = 32'hc13e1809;
    ram_cell[     591] = 32'hd012df8e;
    ram_cell[     592] = 32'ha2da9626;
    ram_cell[     593] = 32'hab45a70c;
    ram_cell[     594] = 32'hbae3f8e4;
    ram_cell[     595] = 32'h1aeea6cb;
    ram_cell[     596] = 32'h319a5c58;
    ram_cell[     597] = 32'hf83ff654;
    ram_cell[     598] = 32'hc1569ba0;
    ram_cell[     599] = 32'hd8565f25;
    ram_cell[     600] = 32'hd3b4b826;
    ram_cell[     601] = 32'h1a13715f;
    ram_cell[     602] = 32'hfb6caa85;
    ram_cell[     603] = 32'ha26e206c;
    ram_cell[     604] = 32'hfed279c7;
    ram_cell[     605] = 32'h73754e84;
    ram_cell[     606] = 32'h50d61735;
    ram_cell[     607] = 32'hdec7c7a3;
    ram_cell[     608] = 32'hbae13736;
    ram_cell[     609] = 32'h0d4ffd15;
    ram_cell[     610] = 32'hab6125d7;
    ram_cell[     611] = 32'h96bb11a6;
    ram_cell[     612] = 32'he2f65f7e;
    ram_cell[     613] = 32'h5730c828;
    ram_cell[     614] = 32'hb01770f8;
    ram_cell[     615] = 32'h71881de4;
    ram_cell[     616] = 32'hb092241d;
    ram_cell[     617] = 32'h1a76c74c;
    ram_cell[     618] = 32'hcdf5e23f;
    ram_cell[     619] = 32'hb8437147;
    ram_cell[     620] = 32'hd595fa9f;
    ram_cell[     621] = 32'hba9ba97f;
    ram_cell[     622] = 32'h2a822f92;
    ram_cell[     623] = 32'hbc6e44ca;
    ram_cell[     624] = 32'hd2b317f8;
    ram_cell[     625] = 32'h348f85a1;
    ram_cell[     626] = 32'h68e5780a;
    ram_cell[     627] = 32'h1badba43;
    ram_cell[     628] = 32'h8f5da2dc;
    ram_cell[     629] = 32'hba0fdfdb;
    ram_cell[     630] = 32'hd2a50a13;
    ram_cell[     631] = 32'h82f0b950;
    ram_cell[     632] = 32'hcf834ae7;
    ram_cell[     633] = 32'h14c76e58;
    ram_cell[     634] = 32'h1ebcc45e;
    ram_cell[     635] = 32'hfa92f136;
    ram_cell[     636] = 32'h35666efb;
    ram_cell[     637] = 32'hda9fda0c;
    ram_cell[     638] = 32'hb92eee76;
    ram_cell[     639] = 32'hc54aa5f5;
    ram_cell[     640] = 32'h07b77c62;
    ram_cell[     641] = 32'he943dd6a;
    ram_cell[     642] = 32'h6f524f8e;
    ram_cell[     643] = 32'hcdb5d7a3;
    ram_cell[     644] = 32'hf502fd54;
    ram_cell[     645] = 32'he66a6fd1;
    ram_cell[     646] = 32'hb5a25c7d;
    ram_cell[     647] = 32'h533d8b58;
    ram_cell[     648] = 32'h162ce617;
    ram_cell[     649] = 32'ha6193ae9;
    ram_cell[     650] = 32'hfa62ebd4;
    ram_cell[     651] = 32'h424e0a4e;
    ram_cell[     652] = 32'h76b0b0b2;
    ram_cell[     653] = 32'hdd5a8f95;
    ram_cell[     654] = 32'h4436ec93;
    ram_cell[     655] = 32'hd2bdbd9d;
    ram_cell[     656] = 32'h22270841;
    ram_cell[     657] = 32'hd7bcbf7e;
    ram_cell[     658] = 32'hc731ddb9;
    ram_cell[     659] = 32'h975f9296;
    ram_cell[     660] = 32'h57fe9c9c;
    ram_cell[     661] = 32'ha0793d0c;
    ram_cell[     662] = 32'h1dbce1bb;
    ram_cell[     663] = 32'h567e99f7;
    ram_cell[     664] = 32'h56403419;
    ram_cell[     665] = 32'h1aa270bc;
    ram_cell[     666] = 32'h2f8663da;
    ram_cell[     667] = 32'hab225480;
    ram_cell[     668] = 32'he5647867;
    ram_cell[     669] = 32'h63e9cf5a;
    ram_cell[     670] = 32'h71124546;
    ram_cell[     671] = 32'h9cd679cf;
    ram_cell[     672] = 32'h2d31824e;
    ram_cell[     673] = 32'h1c3f5949;
    ram_cell[     674] = 32'h23b2fdb7;
    ram_cell[     675] = 32'h90a5e084;
    ram_cell[     676] = 32'h6d1393ed;
    ram_cell[     677] = 32'h0d133c99;
    ram_cell[     678] = 32'h4eb5148d;
    ram_cell[     679] = 32'h4f11e57d;
    ram_cell[     680] = 32'hbe1c636e;
    ram_cell[     681] = 32'ha49fbc7b;
    ram_cell[     682] = 32'ha54ac568;
    ram_cell[     683] = 32'h627ddd5e;
    ram_cell[     684] = 32'h361b4750;
    ram_cell[     685] = 32'h47ddb141;
    ram_cell[     686] = 32'hc5de73d9;
    ram_cell[     687] = 32'h931efd81;
    ram_cell[     688] = 32'h4fcefb61;
    ram_cell[     689] = 32'h41a657e8;
    ram_cell[     690] = 32'hcb9851e8;
    ram_cell[     691] = 32'h0e8d426e;
    ram_cell[     692] = 32'h5180386b;
    ram_cell[     693] = 32'hc675c2d3;
    ram_cell[     694] = 32'h545f3e15;
    ram_cell[     695] = 32'h9ed83f46;
    ram_cell[     696] = 32'h06478526;
    ram_cell[     697] = 32'he0564088;
    ram_cell[     698] = 32'hbdc0283e;
    ram_cell[     699] = 32'h60392ac5;
    ram_cell[     700] = 32'hb42ac129;
    ram_cell[     701] = 32'h8e385f5d;
    ram_cell[     702] = 32'h27837877;
    ram_cell[     703] = 32'hb9536e7f;
    ram_cell[     704] = 32'h4eaa97c1;
    ram_cell[     705] = 32'h14018b0c;
    ram_cell[     706] = 32'hd247ecd1;
    ram_cell[     707] = 32'hefbcebbf;
    ram_cell[     708] = 32'h48544fe7;
    ram_cell[     709] = 32'h3eb2abb8;
    ram_cell[     710] = 32'h32a9ca2b;
    ram_cell[     711] = 32'hebd0ca05;
    ram_cell[     712] = 32'h0714e79f;
    ram_cell[     713] = 32'ha8b2cb2d;
    ram_cell[     714] = 32'hc5d5aa6d;
    ram_cell[     715] = 32'h42d7a332;
    ram_cell[     716] = 32'h5c9976ef;
    ram_cell[     717] = 32'h912fd00a;
    ram_cell[     718] = 32'h4262375a;
    ram_cell[     719] = 32'h4a3fa8ed;
    ram_cell[     720] = 32'hb7bab106;
    ram_cell[     721] = 32'h551b3c02;
    ram_cell[     722] = 32'h13cd61d4;
    ram_cell[     723] = 32'h9e6c8a5e;
    ram_cell[     724] = 32'h4ddeb33f;
    ram_cell[     725] = 32'hcbf2577f;
    ram_cell[     726] = 32'h20386864;
    ram_cell[     727] = 32'h29afe41c;
    ram_cell[     728] = 32'h3fd03666;
    ram_cell[     729] = 32'he74f4215;
    ram_cell[     730] = 32'h2a19717b;
    ram_cell[     731] = 32'h421ac3f9;
    ram_cell[     732] = 32'h3987e96e;
    ram_cell[     733] = 32'hbe04f70c;
    ram_cell[     734] = 32'h108b891a;
    ram_cell[     735] = 32'h2fc01757;
    ram_cell[     736] = 32'h7d634885;
    ram_cell[     737] = 32'h3c56df28;
    ram_cell[     738] = 32'h13b8fd67;
    ram_cell[     739] = 32'h8dca566e;
    ram_cell[     740] = 32'hea209111;
    ram_cell[     741] = 32'h8082b48e;
    ram_cell[     742] = 32'h32859535;
    ram_cell[     743] = 32'h6168eb09;
    ram_cell[     744] = 32'he2e20bf8;
    ram_cell[     745] = 32'hfdd7b8d6;
    ram_cell[     746] = 32'h10b3ab42;
    ram_cell[     747] = 32'h0d1875b6;
    ram_cell[     748] = 32'hb2fb9c52;
    ram_cell[     749] = 32'h11401338;
    ram_cell[     750] = 32'h3cb26424;
    ram_cell[     751] = 32'h868fa150;
    ram_cell[     752] = 32'h4e6f79bb;
    ram_cell[     753] = 32'h643f7916;
    ram_cell[     754] = 32'h1590577b;
    ram_cell[     755] = 32'h4de67588;
    ram_cell[     756] = 32'h64a9788a;
    ram_cell[     757] = 32'h562abb54;
    ram_cell[     758] = 32'ha816d02d;
    ram_cell[     759] = 32'h2b661fa9;
    ram_cell[     760] = 32'hdc61f5f4;
    ram_cell[     761] = 32'hf7d08606;
    ram_cell[     762] = 32'hc89e643f;
    ram_cell[     763] = 32'h09318f1a;
    ram_cell[     764] = 32'h04d8af14;
    ram_cell[     765] = 32'h0bb13a9b;
    ram_cell[     766] = 32'ha011c04c;
    ram_cell[     767] = 32'h034f2273;
end

endmodule

